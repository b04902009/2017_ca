module Instruction_Memory(
    addr_i, 
    instr_o
);

// Interface
input   [31:0]      addr_i;
output  [31:0]      instr_o;

// Instruction memory
reg     [31:0]     memory  [0:255]; // Declaration of 256 32-bit registers

assign  instr_o = memory[addr_i>>2];  
// always @(*) begin
// 	$display("Instruction_Memory-instr: %b", instr_o);
// end

endmodule
